module main;
    initial
        begin
            $display("Learning Verilog");
            $finish;
        end
endmodule
